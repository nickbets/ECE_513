* First line should be ignored

* Voltage Sources
V1 n_A 0 5
V2 3 n_2 0.3
V3 n_X 6 1.5

* Current Sources
I1 4 n_Y 2e-3
I2 n_B 6 1e-3

* Resistors
R1 1 n_A 1.8
R2 1 n_2 1.2
R3 n_A n_2 75
R4 n_2 n_X 0.2
R5 n_2 6 2.5
R6 3 n_Y 0.15
R7 n_Y 0 5e2
R8 n_X 0 15
R9 3 n_4_4 10
R10 nodeC n_B 8.3

* Capacitors
C1 1 n_2 4e-6
C2 3 n_X 2e-6
C3 n_A n_Y 5e-6

* Inductors
L1 n_2 nodeZ 7e-3
L2 nodeZ 7 12e-3
L3 n_X 0 3e-3

* Diodes with Optional Area Parameter
D1 4 n_A DModel area=1.2
D2 n_B 0 DModel

* MOSFET Transistors
M1 n_2 3 n_4_4 0 NMOS L=2e-6 W=8e-6
M2 nodeC n_A 4 0 PMOS L=1e-6 W=15e-6

* BJT Transistors with Optional Area Parameter
Q1 n_X n_2 0 QModel area=1.5
Q2 n_4_4 n_Y 0 PModel

*** .MODEL command is optional since it will not be used in this course ***
*.MODEL DModel D IS=1e-14
*.MODEL NMOS NMOS LEVEL=1 VTO=0.7 KP=120u
*.MODEL PMOS PMOS LEVEL=1 VTO=-0.8 KP=90u
*.MODEL QModel NPN IS=1e-15 BF=150
*.MODEL PModel PNP IS=1e-15 BF=100

* usually we define the EOF with .END but it's optional
*.END